module top_module (
	input clk,
	input d,
	input ar,
	output logic q
);


endmodule
